`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "apb_interface.sv"
`include "apb_sequence_items.sv"
`include "apb_sequence.sv"
`include "apb_sequencer.sv"
`include "apb_driver.sv"
`include "apb_monitor.sv"
`include "apb_scorboard.sv"
`include "apb_agent.sv"
`include "apb_coverage.sv"
`include "apb_environment.sv"
`include "apb_test.sv"


